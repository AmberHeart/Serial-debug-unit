// `timescale 1ns / 1ps

// module uart_rx(
//     input clk,//9600*16  HZ
//     input rstn,
//     input rxd,
//     input rdy_rx,//1 means ready to accept new data, 0 otherwise.pulse signal
//     output reg [7:0] d_rx,
//     output reg vld_rx   //1 indicates that data has been received and is waiting for other modules to take it away
// );

// // parameter TICKS_PER_BIT = 10416; // assuming 100 MHz clock frequency
// reg [15:0] CNT;
// // reg[3:0] fr_div;//分频器
// reg [3:0] CNTb;
// wire process;//表示是否正在接收数据，1表示正在接受
// assign flg=process;
// CNTc cntc(
//     /*
//     input clk,
//     input rstn,
//     input rxd,
//     input vld_rx,
//     output reg process
//     */
//     .clk(clk),
//     .rstn(rstn),
//     .rxd(rxd),
//     .vld_rx(vld_rx),//vld_rx=1--->process=0
//     .process(process)
// );
// reg edg_up,tmp;//取process上升沿
// always @(posedge clk) begin
//     tmp<=process;
//     if(process&&!tmp)begin
//         edg_up<=1;
//     end else begin
//         edg_up<=0;
//     end
// end
// always @(posedge clk) begin
//     if(rstn||edg_up||rdy_rx)begin
//         d_rx<=0;
//         CNT<=0;
//     end
//     if(process) begin
//         if(CNT==8)begin//取样中点
//             CNT<=0;
//             d_rx<={rxd,d_rx[7:1]};
//         end else begin
//             CNT<=CNT+1;
//         end
//     end
// end
// always @(posedge clk) begin
//     if(rstn||edg_up||rdy_rx)begin
//         CNTb<=0;
//         vld_rx<=0;
//     end else if(process)begin
//         if(CNT==0)begin//取样中数据还未被接受
//             CNTb<=CNTb+1;
//         end
//         if(CNTb==8)begin
//             vld_rx<=1;
//             CNTb<=0;
//         end else begin
//             vld_rx<=0;
//         end
//     end 
// end
// endmodule   
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/03/20 14:51:12
// Design Name: 
// Module Name: RX
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module RX(
    input clk,//16*9600Hz
    input rstn,
    input rxd,//urat signal
    output reg vld_rx,//1 indicates that data has been received and is waiting for other modules to take it away
    input rdy_rx,//1 means ready to accept new data, 0 otherwise.
    output [7:0] d_rx
    );
    // //100MHZ change to 16*9600 HZ 
    wire div_clk = clk;
    /*DIV_RX_CLK div_rx_clk(
        .clk(clk),
        .rstn(rstn),
        .div_clk(div_clk)
    );*/
    //Shift Input Register
    wire SIR_saved;
    wire [8:0] SIR;
    SIR sir(
        .clk(div_clk),
        .rstn(rstn),
        .rxd(rxd),
        .SIR_saved(SIR_saved),
        .SIR(SIR)
    );
    reg [7:0] DIR;
    always@(posedge clk)
    begin
        if(vld_rx == 0)
        begin
            if(SIR_saved == 1)
            begin
                vld_rx <= 1;
                DIR <= SIR[7:0];
            end
            else //no data 
                DIR <= 8'h00;
        end
        else
        begin
            if(rdy_rx == 1)
                vld_rx <= 0;
            else
                vld_rx <= vld_rx;
        end
    end
    assign d_rx = DIR;
endmodule
