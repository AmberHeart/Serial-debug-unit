`timescale 1ns / 1ps
module DCP_G(
    input clk,
    input rstn,
    input [7:0] sel_mode,
    input [7:0] CMD_G,
    output reg finish_G,
    input [31:0] pc_chk,
    input [31:0] B_1,
    input [31:0] B_2,
    input [31:0] din_rx,
    input flag_rx,
    input ack_rx,
    output reg req_rx_G,
    output type_rx_G,
    output reg clk_cpu_G,

    input [31:0] IMM, // immed
    input [31:0] pc, // curren
    input [31:0] npc, //next p
    input [31:0] IR, // instru
    input [31:0] CTL, // contr
    input [31:0] A, // registe
    input [31:0] B, // registe
    input [31:0] Y, // ALU res
    input [31:0] MDR, // memor
    input ack_tx,
    output reg req_tx_G,
    output reg type_tx_G,
    output reg [31:0] dout_G
);

assign type_rx_G = 0;
    // always@(*) begin
    //     if(pc_chk == B_1 || pc_chk == B_2 || din_rx == 8'h48) begin
    //         finish_G=1;
    //         clk_cpu_G_G = 0;
    //     end
    //     else begin
    //         finish_G=0;
    //         clk_cpu_G_G = clk;
    //     end
    // end
    // always@(posedge clk or negedge rstn) begin
    //     if(~rstn) begin
    //         req_rx_G<=0;
    //     end
    //     else begin
    //         if (sel_mode == CMD_G) begin
    //             if(~ack_rx) begin
    //                 req_rx_G<=1;
    //             end
    //             else begin
    //                 req_rx_G<=0;
    //             end
    //         end
    //     end
    
    // end
        parameter [4:0]
    INIT = 5'b00000,
    CLK_ON = 5'b10100,
    PRINT_NPC = 5'b00001,
    PRINT_NPC_DATA = 5'b00010,
    PRINT_PC = 5'b00011,
    PRINT_PC_DATA = 5'b00100,
    PRINT_IR = 5'b00101,
    PRINT_IR_DATA = 5'b00110,
    PRINT_CTL = 5'b00111,
    PRINT_CTL_DATA = 5'b01000,
    PRINT_A = 5'b01001,
    PRINT_A_DATA = 5'b01010,
    PRINT_B = 5'b01011,
    PRINT_B_DATA = 5'b01100,
    PRINT_IMM = 5'b01101,
    PRINT_IMM_DATA = 5'b01110,
    PRINT_Y = 5'b01111,
    PRINT_Y_DATA = 5'b10000,
    PRINT_MDR = 5'b10001,
    PRINT_MDR_DATA = 5'b10010,
    FINISH = 5'b10011;
    reg [4:0] CS=INIT, NS=INIT;
    //PRINT
    reg [2:0] count_NPC=0;
    reg [2:0] count_PC=0;
    reg [2:0] count_IR=0;
    reg [2:0] count_CTL=0;
    reg [2:0] count_A=0;
    reg [2:0] count_B=0;
    reg [2:0] count_IMM=0;
    reg [2:0] count_Y=0;
    reg [2:0] count_MDR=0;
    reg count_FINISH =0;
    wire we;
    assign we = (sel_mode == CMD_G);
    always @(posedge clk or negedge rstn) begin
        if(~rstn) begin
            CS<=INIT;
            finish_G<=0;
            count_NPC<=0;
            count_PC<=0;
            count_IR<=0;
            count_CTL<=0;
            count_A<=0;
            count_B<=0;
            count_IMM<=0;
            count_Y<=0;
            count_MDR<=0;
            //req_rx_P<=0;
            req_tx_G<=0;
        end
        else begin 
            CS<=NS;
            case(CS)
                INIT: begin
                    finish_G<=0;
                    count_NPC<=0;
                    count_PC<=0;
                    count_IR<=0;
                    count_CTL<=0;
                    count_A<=0;
                    count_B<=0;
                    count_IMM<=0;
                    count_Y<=0;
                    count_MDR<=0;
                    //req_rx_P<=0;
                    count_FINISH <=0;
                    clk_cpu_G <=0;
                end
                CLK_ON: begin
                    clk_cpu_G <=~clk_cpu_G;
                    if (~ack_rx) begin
                        req_rx_G <= 1;
                    end
                    else begin
                        req_rx_G <= 0;
                        
                    end
                end
                
                PRINT_NPC: begin
                    if(count_NPC < 3) begin
                        if(ack_tx) begin
                            count_NPC <=count_NPC + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_NPC <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_NPC_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                PRINT_PC: begin
                    if(count_PC < 2) begin
                        if(ack_tx) begin
                            count_PC <=count_PC + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_PC <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_PC_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                PRINT_IR: begin
                    if(count_IR < 2) begin
                        if(ack_tx) begin
                            count_IR <=count_IR + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_IR <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_IR_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                PRINT_CTL: begin
                    if(count_CTL < 3) begin
                        if(ack_tx) begin
                            count_CTL <=count_CTL + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_CTL <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_CTL_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                PRINT_A: begin
                    if(count_A < 1) begin
                        if(ack_tx) begin
                            count_A <=count_A + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_A <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_A_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                PRINT_B: begin
                    if(count_B < 1) begin
                        if(ack_tx) begin
                            count_B <=count_B + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_B <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_B_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                PRINT_IMM: begin
                    if(count_IMM < 3) begin
                        if(ack_tx) begin
                            count_IMM <=count_IMM + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_IMM <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_IMM_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                PRINT_Y: begin
                    if(count_Y < 1) begin
                        if(ack_tx) begin
                            count_Y <=count_Y + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_Y <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_Y_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                PRINT_MDR: begin
                    if(count_MDR < 3) begin
                        if(ack_tx) begin
                            count_MDR <=count_MDR + 1;
                            req_tx_G<=0;
                        end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_MDR <= 0;
                            req_tx_G <= 0;
                        end
                        else req_tx_G <= 1;
                    end
                end
                PRINT_MDR_DATA: begin
                    if(ack_tx) begin
                        req_tx_G <= 0;
                    end
                    else req_tx_G <= 1;
                end
                FINISH: begin
                    if(count_FINISH == 0) begin
                        if(ack_tx) begin
                            count_FINISH <= 1;
                            req_tx_G<=0;
                    end
                        else req_tx_G<=1;
                    end
                    else begin
                        if (ack_tx) begin
                            count_FINISH <= 0;
                            req_tx_G <= 0;
                            finish_G <= 1;
                        end
                        else req_tx_G <= 1;
                    end
                end
                default begin
                            CS<=INIT;
                            finish_G<=0;
                            count_NPC<=0;
                            count_PC<=0;
                            count_IR<=0;
                            count_CTL<=0;
                            count_A<=0;
                            count_B<=0;
                            count_IMM<=0;
                            count_Y<=0;
                            count_MDR<=0;
                            //req_rx_P<=0;
                            req_tx_G<=0;
                end
            endcase
        end
    end
    always @(*) begin
        type_tx_G = 0;
        dout_G = 0;
        NS = INIT;
        if(~we) NS =INIT;
        
        else case (CS)
            INIT: begin
                if(we) NS = CLK_ON;
                else NS = INIT;
            end
            CLK_ON: begin
                if(din_rx == 32'h48 || pc_chk == B_1 || pc_chk == B_2) begin
                    NS = PRINT_NPC;
                end
                else NS=CLK_ON;
                
            end
            
            PRINT_NPC: begin //ASCII_NPC <= 32'h4E50433D;//NPC=
                if(count_NPC == 0) begin
                     NS = PRINT_NPC;
                     type_tx_G = 0;
                     dout_G=32'h4E;
                end
                else if(count_NPC == 1) begin
                    NS = PRINT_NPC;
                    type_tx_G = 0;
                    dout_G=32'h50;
                end
                else if(count_NPC == 2) begin
                    NS = PRINT_NPC;
                    type_tx_G = 0;
                    dout_G=32'h43;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_NPC_DATA;
                    end
                    else NS = PRINT_NPC;
                end
            end
            PRINT_NPC_DATA: begin
                type_tx_G = 1;
                dout_G = npc;
                if(~ack_tx) NS = PRINT_NPC_DATA;
                else NS = PRINT_PC;
            end
            PRINT_PC: begin //ASCII_PC <= 32'h50433D;//PC=
                if(count_PC == 0) begin
                     NS = PRINT_PC;
                     type_tx_G = 0;
                     dout_G=32'h50;
                end
                else if(count_PC == 1) begin
                    NS = PRINT_PC;
                    type_tx_G = 0;
                    dout_G=32'h43;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_PC_DATA;
                    end
                    else NS = PRINT_PC;
                end
            end
            PRINT_PC_DATA: begin
                type_tx_G = 1;
                dout_G = pc;
                if(~ack_tx) NS = PRINT_PC_DATA;
                else NS = PRINT_IR;
            end
            PRINT_IR: begin //ASCII_IR <= 32'h49523D;//IR=
                if(count_IR == 0) begin
                     NS = PRINT_IR;
                     type_tx_G = 0;
                     dout_G=32'h49;
                end
                else if(count_IR == 1) begin
                    NS = PRINT_IR;
                    type_tx_G = 0;
                    dout_G=32'h52;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_IR_DATA;
                    end
                    else NS = PRINT_IR;
                end
            end
            PRINT_IR_DATA: begin
                type_tx_G = 1;
                dout_G = IR;
                if(~ack_tx) NS = PRINT_IR_DATA;
                else NS = PRINT_CTL;
            end
            PRINT_CTL: begin //ASCII_CTL <= 32'h43544C3D;
                if(count_CTL == 0) begin
                     NS = PRINT_CTL;
                     type_tx_G = 0;
                     dout_G=32'h43;
                end
                else if(count_CTL == 1) begin
                    NS = PRINT_CTL;
                    type_tx_G = 0;
                    dout_G=32'h54;
                end
                else if(count_CTL == 2) begin
                    NS = PRINT_CTL;
                    type_tx_G = 0;
                    dout_G=32'h4C;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_CTL_DATA;
                    end
                    else NS = PRINT_CTL;
                end
            end
            PRINT_CTL_DATA: begin
                type_tx_G = 1;
                dout_G = CTL;
                if(~ack_tx) NS = PRINT_CTL_DATA;
                else NS = PRINT_A;
            end
            PRINT_A: begin //ASCII_A <= 32'h413D;//A=
                if(count_A == 0) begin
                     NS = PRINT_A;
                     type_tx_G = 0;
                     dout_G=32'h41;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_A_DATA;
                    end
                    else NS = PRINT_A;
                end
            end
            PRINT_A_DATA: begin
                type_tx_G = 1;
                dout_G = A;
                if(~ack_tx) NS = PRINT_A_DATA;
                else NS = PRINT_B;
            end
            PRINT_B: begin //ASCII_B <= 32'h423D;//B=
                if(count_B == 0) begin
                     NS = PRINT_B;
                     type_tx_G = 0;
                     dout_G=32'h42;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_B_DATA;
                    end
                    else NS = PRINT_B;
                end
            end
            PRINT_B_DATA: begin
                type_tx_G = 1;
                dout_G = B;
                if(~ack_tx) NS = PRINT_B_DATA;
                else NS = PRINT_IMM;
            end
            PRINT_IMM: begin //ASCII_IMM <= 32'h494D4D3D;//IMM=
                if(count_IMM == 0) begin
                     NS = PRINT_IMM;
                     type_tx_G = 0;
                     dout_G=32'h49;
                end
                else if(count_IMM == 1) begin
                    NS = PRINT_IMM;
                    type_tx_G = 0;
                    dout_G=32'h4D;
                end
                else if(count_IMM == 2) begin
                    NS = PRINT_IMM;
                    type_tx_G = 0;
                    dout_G=32'h4D;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_IMM_DATA;
                    end
                    else NS = PRINT_IMM;
                end
            end
            PRINT_IMM_DATA: begin
                type_tx_G = 1;
                dout_G = IMM;
                if(~ack_tx) NS = PRINT_IMM_DATA;
                else NS = PRINT_Y;
            end
            PRINT_Y: begin //ASCII_Y <= 32'h593D;//Y=
                if(count_Y == 0) begin
                     NS = PRINT_Y;
                     type_tx_G = 0;
                     dout_G=32'h59;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_Y_DATA;
                    end
                    else NS = PRINT_Y;
                end
            end
            PRINT_Y_DATA: begin
                type_tx_G = 1;
                dout_G = Y;
                if(~ack_tx) NS = PRINT_Y_DATA;
                else NS = PRINT_MDR;
            end
            PRINT_MDR: begin //ASCII_MDR <= 32'h4D44523D;//MDR=
                if(count_MDR == 0) begin
                     NS = PRINT_MDR;
                     type_tx_G = 0;
                     dout_G=32'h4D;
                end
                else if(count_MDR == 1) begin
                    NS = PRINT_MDR;
                    type_tx_G = 0;
                    dout_G=32'h44;
                end
                else if(count_MDR == 2) begin
                    NS = PRINT_MDR;
                    type_tx_G = 0;
                    dout_G=32'h52;
                end
                else  begin
                    type_tx_G = 0;
                    dout_G=32'h3D;
                    if(ack_tx) begin
                        NS=PRINT_MDR_DATA;
                    end
                    else NS = PRINT_MDR;
                end
            end
            PRINT_MDR_DATA: begin
                type_tx_G = 1;
                dout_G = MDR;
                if(~ack_tx) NS = PRINT_MDR_DATA;
                else NS = FINISH;
            end
            FINISH: begin
                if (count_FINISH == 0) begin
                    type_tx_G = 0;
                    dout_G = 32'h0d;
                    NS = FINISH;
                end
                else begin
                    type_tx_G = 0;
                    dout_G = 32'h0a;
                    if (ack_tx) begin
                        NS = INIT;
                        
                    end
                    else NS = FINISH;
                end
            end


            endcase
    end
    //assign cs=CS;
endmodule