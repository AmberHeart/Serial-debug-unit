`timescale 1ps/1ps

module test();
    input reg [7:0] a;
    output    [7:0] b;
    assign b = a;
endmodule
